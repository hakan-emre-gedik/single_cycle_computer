module memory_128x8bit(
	data_out, 
	data_in, 
	address_in, 
	we
); 
	output reg [31:0] data_out; // input and output should have 32-bit length. 	
	input [31:0] data_in; 
	input [31:0] address_in; 
	input we; 

	reg [31:0] mem[127:0]; 
	
	always @(*) begin 
		if (we) begin 
			mem[address_in] <= data_in; 
		end 
		data_out <= mem[address_in]; 
	end 

endmodule 